SIMPLPARAEQ (TINA Netlist Editor format)
**************************************
**  This file was created by TINA   **
**         www.tina.com             ** 
**      (c) DesignSoft, Inc.        **          
**     www.designsoftware.com       **
**************************************
.LIB "<TINADIR>\EXAMPLES\SPICE\TSPICE.LIB"
.LIB "<TINADIR>\SPICELIB\Operational Amplifiers.LIB"
.TEMP 27
.AC DEC 33 20 20K
.TRAN 2N 1U
.DC LIN Vin 0 1 10M

.PROBE V([Vout])

Vnegdc      0 3 15
Vposdc      2 0 15
Vin         13 0 DC 0 AC 1 0
+ PULSE ( 0 1 0  0  0  1e19 1e20 )
XU4         0 1 2 3 4 OPA1612_0
XU5         0 5 2 3 Vout OPA1612_0
XU1         0 7 2 3 8 OPA1612_0
XU2         0 9 2 3 10 OPA1612_0
XU3         0 11 2 3 12 OPA1612_0
C2          11 12 10N 
C1          9 10 10N 
XPboostcut   13 Vout 14  PotMeter PARAMS: Res=10K Percent=10M
Rq2         1 10 1K 
R7          4 1 1K 
R6          4 7 1K 
Rq1         14 7 1K 
R3          12 7 1K 
R2          7 8 1K 
Rfr1        8 9 15K 
Rfr2        10 11 15K 
R5          5 Vout 1K 
R4          13 5 1K 
Rbcmax      10 5 1K 


.LIB "<TINADIR>\SPICELIB\Operational Amplifiers.LIB"
*$
* OPA1612
*$
*****************************************************************************
* (C) COPYRIGHT 2011 TEXAS INSTRUMENTS INCORPORATED. ALL RIGHTS RESERVED.                                            
*****************************************************************************
** THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.
** TI AND ITS LICENSORS AND SUPPLIERS MAKE NO WARRANTIES, EITHER EXPRESSED
** OR IMPLIED, WITH RESPECT TO THIS MODEL, INCLUDING THE WARRANTIES OF 
** MERCHANTABILITY OR FITNESS FOR A PARTICULAR PURPOSE.  THE MODEL IS
** PROVIDED SOLELY ON AN "AS IS" BASIS.  THE ENTIRE RISK AS TO ITS QUALITY
** AND PERFORMANCE IS WITH THE CUSTOMER.
*****************************************************************************
*
* THIS MODEL IS SUBJECT TO CHANGE WITHOUT NOTICE. TEXAS INSTRUMENTS
* INCORPORATED IS NOT RESPONSIBLE FOR UPDATING THIS MODEL.
*
*****************************************************************************
*
** RELEASED BY: ANALOG ELAB DESIGN CENTER, TEXAS INSTRUMENTS INC.
* PART: OPA1612
* DATE: 13JUN2011
* MODEL TYPE: ALL IN ONE
* SIMULATOR: TINA
* SIMULATOR VERSION: 9.1.30.94 SF-TI
* EVM ORDER NUMBER: N/A
* EVM USERS GUIDE: N/A
* DATASHEET: SBOS450A�JULY 2009�REVISED AUGUST 2009
*
* MODEL VERSION: 1.0
*
*****************************************************************************
* 
* UPDATES:
*
* VERSION 1.0 : 
* RELEASE TO WEB
*
*****************************************************************************
* COMMENTS:
*
* MODEL FEATURES INCLUDE OUTPUT SWING, OUTPUT CURRENT THROUGH
* THE SUPPLY RAILS, RAIL-TO-RAIL OUTPUT STAGE, OUTPUT CURRENT
* LIMIT, OPEN LOOP GAIN AND PHASE WITH RL AND CL EFFECTS,
* SLEW RATE WITH TEMPERATURE EFFECTS, SETTLING TIME TO 0.01 %,
* OVERLOAD RECOVERY TIME, COMMON MODE REJECTION WITH FREQUENCY
* EFFECTS, OUTPUT IMPEDANCE, POWER SUPPLY REJECTION WITH
* FREQUENCY EFFECTS, INPUT VOLTAGE NOISE WITH 1/F AND FEATURE
* AT 20 MEGAHERTZ, INPUT CURRENT NOISE WITH 1/F, INPUT BIAS
* CURRENT, INPUT IMPEDANCE, INPUT COMMON MODE RANGE, INPUT
* OFFSET VOLTAGE WITH TEMPERATURE EFFECTS, AND QUIESCENT
* CURRENT VS VOLTAGE AND TEMPERATURE. MODEL INCLUDES INPUT
* PROTECTION DIODES.
* MODEL DOES NOT INCLUDE SHUTDOWN.
* THIS MODEL IS ALSO APPLICABLE TO OPA1611.
*
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  3   2   7  4  6
*****************************************************************************
.SUBCKT OPA1612_0  3 2 7 4 6
D17 9 0 DIN
D18 10 0 DIN
I14 0 9 0.1E-3
I15 0 10 0.1E-3
D19 11 0 DVN
D20 12 0 DVN
I16 0 11 0.1E-3
I17 0 12 0.1E-3
E15 13 14 11 12 4.23E-2
G5 15 13 9 10 1.1E-4
E16 16 0 17 0 1
E17 18 0 19 0 1
E18 20 0 21 0 1
R56 16 22 1E6
R57 18 23 1E6
R58 20 24 1E4
R59 0 22 10
R60 0 23 10
R61 0 24 7
E19 25 26 27 0 0.1
R62 28 21 1E3
R63 21 29 1E3
C15 16 22 1E-12
C16 18 23 1E-12
C17 20 24 1E-9
E20 30 25 23 0 -1E-3
E21 31 30 22 0 1E-3
R64 0 32 1E12
G12 15 13 33 0 1.45E-14
R136 0 33 10E3
R137 0 33 10E3
R138 26 25 1E9
R139 25 30 1E9
R140 30 31 1E9
E74 29 0 15 0 1
E75 28 0 13 0 1
C23 15 13 0.05E-12
E77 26 3 34 0 1.98E-4
R146 26 3 1E9
R147 0 32 1E12
Q41 35 36 19 QLN
R148 36 37 1E3
R149 38 39 1E3
R150 40 17 5
R151 19 41 5
R153 42 43 850
R154 44 17 5
R155 19 45 5
D22 46 7 DD
D23 4 46 DD
E58 19 0 4 0 1
E79 17 0 7 0 1
R156 4 7 1.1E9
E60 47 19 17 19 0.5
D24 48 17 DD
D25 19 49 DD
R157 50 51 100
R158 52 53 100
G14 42 47 54 47 0.1E-3
R159 47 42 5.3E6
C24 43 55 5P
C25 46 0 0.5E-12
D26 53 35 DD
D27 56 51 DD
Q42 56 39 17 QLP
R160 46 57 1
R161 58 46 1
E71 59 47 60 61 1
R162 59 54 1E4
C26 54 47 0.02P
G15 62 47 42 47 -1E-3
G16 47 63 42 47 1E-3
G17 47 64 65 19 1E-3
G18 66 47 17 67 1E-3
D28 66 62 DD
D29 63 64 DD
R163 62 66 100E6
R164 64 63 100E6
R165 66 17 1E3
R166 19 64 1E3
R167 63 47 1E6
R168 64 47 1E6
R169 47 66 1E6
R170 47 62 1E6
G19 7 4 68 0 3.5E-3
R171 47 54 1E9
R172 50 17 1E9
R173 19 52 1E9
G20 67 65 32 0 1E-3
L2 46 6 0.4E-9
R175 46 6 400
R176 67 17 1E8
R177 19 65 1E8
R178 41 53 1E8
R179 40 51 1E8
R180 0 32 1E9
E84 17 38 17 40 5
E85 37 19 41 19 3
E24 55 0 46 0 1
R219 42 55 1.8E9
I30 0 69 1E-3
D46 69 0 DD
R278 0 69 10E6
V27 69 34 0.65
R279 0 34 10E6
Q52 57 51 40 QOP
Q53 58 53 41 QON
Q54 65 65 45 QON
Q55 67 67 44 QOP
E144 17 50 17 66 1
E145 52 19 64 19 1
Q56 70 15 71 QIN
Q57 72 13 73 QIN
Q58 61 74 70 QIN
Q59 60 75 72 QIN
Q60 74 74 76 QIP
Q61 15 74 76 QIP
Q62 75 75 76 QIP
Q63 13 75 76 QIP
R280 61 77 1200
R281 60 77 1200
R282 78 71 4
R283 78 73 4
Q64 78 79 80 QTN
C108 61 81 1E-15
R284 81 55 600
I33 0 82 1E-3
D49 82 0 DD
R287 0 82 10E6
V30 82 83 1.2301
R288 0 83 10E6
E50 84 0 83 0 -1.75
R289 0 84 10E6
R290 85 84 10E6
M3 85 86 0 0 NEN L=2U W=1000U
G22 80 79 85 0 12E-6
V32 87 0 1
R291 87 86 1E6
M4 86 32 0 0 NEN L=2U W=100U
C109 61 60 4.75E-12
V34 77 76 1
E51 42 49 47 19 0.7
E52 48 42 17 47 0.7
G23 7 0 57 46 1
G24 4 0 46 58 -1
V35 17 8 1
M45 88 89 90 90 NEN L=3U W=3000U
R293 90 91 1E4
R294 88 17 1E6
V36 17 90 1
C110 17 8 1E-12
E53 32 0 92 90 1
V37 88 92 1.111E-6
R295 90 92 1E12
R296 8 17 1E6
C111 91 90 3E-15
C112 17 88 3E-15
M50 93 94 90 90 NEN L=3U W=300U
M51 89 93 90 90 NEN L=3U W=300U
R297 93 17 1E4
R298 89 17 1E4
C113 17 93 55E-12
C114 17 89 150E-12
E54 95 42 32 0 30
E55 96 47 32 0 -30
V38 97 96 15
V39 98 95 -15
R300 95 0 1E12
R301 96 0 1E12
M52 47 98 42 99 PSW L=1.5U W=150U
M53 42 97 47 100 NSW L=1.5U W=150U
R302 99 0 1E12
R303 100 0 1E12
M54 91 8 17 17 PEN L=6U W=60U
E56 101 90 91 90 -1
R304 90 101 10E6
R305 90 101 10E6
V40 94 101 1
R306 90 94 10E6
E57 102 0 24 0 1
R307 102 27 1E4
R308 0 27 7
C115 102 27 1E-9
M55 103 104 4 4 NEN L=2U W=1000U
R309 103 7 160E3
E78 104 4 32 0 3
V41 80 19 1.23
V42 17 76 0.48
R310 105 13 100
M56 68 106 0 0 NEN L=2U W=10M
R311 68 84 850E3
E70 107 0 32 0 -1
R312 0 107 10E6
R313 0 107 10E6
V43 106 107 1
R314 0 106 10E6
G25 7 4 32 0 -0.85E-3
G26 7 4 108 0 -4E-5
E61 109 0 7 4 1
M57 108 106 0 0 NEN L=2U W=10M
R315 108 109 75E3
E62 2 14 110 0 0.93
R317 0 110 1E3
C116 110 0 2.4E-12
L5 0 110 40E-6
R318 14 2 1E9
C117 0 15 6E-12
C118 13 0 6E-12
V44 31 15 -29E-6
J2 105 15 105 JC
J3 15 105 15 JC
.MODEL JC NJF IS=1E-18
.MODEL QON NPN RC=5
.MODEL QOP PNP RC=5
.MODEL DD D
.MODEL QIN NPN BF=235
.MODEL QIP PNP BF=235
.MODEL QTN NPN
.MODEL DVN D KF=2.5E-15
.MODEL DIN D KF=1E-15
.MODEL QLN NPN
.MODEL QLP PNP
.MODEL NEN NMOS KP=200U VTO=0.5 IS=1E-18
.MODEL PEN PMOS KP=200U VTO=-0.7 IS=1E-18
.MODEL PSW PMOS KP=200U VTO=-7.5 IS=1E-18
.MODEL NSW NMOS KP=200U VTO=7.5 IS=1E-18
.ENDS OPA1612_0 


.END
